-- 32*32 register file
